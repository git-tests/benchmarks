--=============================================================================
--! @file fmcTLU_pkg_body.vhd
--=============================================================================
---
--! @brief VHDL Package Body fmc_mTLU_lib.fmcTLU
--
--! @author  phdgc
--! @date  16:45:08 11/08/12         
--
-- using Mentor Graphics HDL Designer(TM) 2010.3 (Build 21)
--
PACKAGE BODY fmcTLU IS
END fmcTLU;
