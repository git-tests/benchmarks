`timescale 1ns/1ns

module pc036a_fmc_lpc_connector (fmc_prsnt_m2c_l, fmc_pwr_good_flash_rst_b, fmc_tdo, dp0_c2m, \dp0_c2m* , dp0_m2c, \dp0_m2c* , 
    fmc_clk0_m2c, \fmc_clk0_m2c* , fmc_clk1_m2c, \fmc_clk1_m2c* , fmc_la, \fmc_la* , iic_sda_main, fmc_tck_buf, 
    fmc_tms_buf, fpga_tdo, ga0, ga1, gbtclk0_m2c, \gbtclk0_m2c* , gnd, iic_scl_main, p2v5, p3v3, p12v, trst_l, 
    vref_a_m2c );
// generated by  HDL Direct 16.3-S013 (v16-3-85Y) 7/19/2010
// on Fri Mar  4 11:47:41 2011
// from fmc_tlu_v1_lib/PC036A_FMC_LPC_CONNECTOR/sch_1

  output  fmc_prsnt_m2c_l;
  output  fmc_pwr_good_flash_rst_b;
  output  fmc_tdo;
  inout  dp0_c2m;
  inout  \dp0_c2m* ;
  inout  dp0_m2c;
  inout  \dp0_m2c* ;
  inout  fmc_clk0_m2c;
  inout  \fmc_clk0_m2c* ;
  inout  fmc_clk1_m2c;
  inout  \fmc_clk1_m2c* ;
  inout [33:0] fmc_la;
  inout [33:0] \fmc_la* ;
  inout  iic_sda_main;
  input  fmc_tck_buf;
  input  fmc_tms_buf;
  input  fpga_tdo;
  input  ga0;
  input  ga1;
  input  gbtclk0_m2c;
  input  \gbtclk0_m2c* ;
  input  gnd;
  input  iic_scl_main;
  input  p2v5;
  input  p3v3;
  input  p12v;
  input  trst_l;
  input  vref_a_m2c;

  wire  page1_dp0_c2m;
  wire  \page1_dp0_c2m* ;
  wire  page1_dp0_m2c;
  wire  \page1_dp0_m2c* ;
  wire  page1_fmc_clk0_m2c;
  wire  \page1_fmc_clk0_m2c* ;
  wire  page1_fmc_clk1_m2c;
  wire  \page1_fmc_clk1_m2c* ;
  wire [33:0] page1_fmc_la;
  wire [33:0] \page1_fmc_la* ;
  wire  page1_fmc_prsnt_m2c_l;
  wire  page1_fmc_pwr_good_flash_rst_b;
  wire  page1_fmc_tck_buf;
  wire  page1_fmc_tdo;
  wire  page1_fmc_tms_buf;
  wire  page1_fpga_tdo;
  wire  page1_ga0;
  wire  page1_ga1;
  wire  page1_gbtclk0_m2c;
  wire  \page1_gbtclk0_m2c* ;
  wire  page1_gnd;
  wire  page1_iic_scl_main;
  wire  page1_iic_sda_main;
  wire  page1_p12v;
  wire  page1_p2v5;
  wire  page1_p3v3;
  wire  page1_trst_l;
  wire  page1_vref_a_m2c;

  assign page1_dp0_c2m = dp0_c2m;
  assign \page1_dp0_c2m*  = \dp0_c2m* ;
  assign page1_dp0_m2c = dp0_m2c;
  assign \page1_dp0_m2c*  = \dp0_m2c* ;
  assign page1_fmc_clk0_m2c = fmc_clk0_m2c;
  assign \page1_fmc_clk0_m2c*  = \fmc_clk0_m2c* ;
  assign page1_fmc_clk1_m2c = fmc_clk1_m2c;
  assign \page1_fmc_clk1_m2c*  = \fmc_clk1_m2c* ;
  assign page1_fmc_la[5:5] = fmc_la[5:5];
  assign page1_fmc_la[9:9] = fmc_la[9:9];
  assign page1_fmc_la[13:13] = fmc_la[13:13];
  assign page1_fmc_la[33:33] = fmc_la[33:33];
  assign page1_fmc_la[31:31] = fmc_la[31:31];
  assign page1_fmc_la[29:29] = fmc_la[29:29];
  assign page1_fmc_la[0:0] = fmc_la[0:0];
  assign page1_fmc_la[6:6] = fmc_la[6:6];
  assign page1_fmc_la[10:10] = fmc_la[10:10];
  assign page1_fmc_la[18:18] = fmc_la[18:18];
  assign page1_fmc_la[27:27] = fmc_la[27:27];
  assign page1_fmc_la[14:14] = fmc_la[14:14];
  assign page1_fmc_la[26:26] = fmc_la[26:26];
  assign page1_fmc_la[32:32] = fmc_la[32:32];
  assign page1_fmc_la[28:28] = fmc_la[28:28];
  assign page1_fmc_la[30:30] = fmc_la[30:30];
  assign page1_fmc_la[2:2] = fmc_la[2:2];
  assign page1_fmc_la[19:19] = fmc_la[19:19];
  assign page1_fmc_la[24:24] = fmc_la[24:24];
  assign page1_fmc_la[21:21] = fmc_la[21:21];
  assign page1_fmc_la[3:3] = fmc_la[3:3];
  assign page1_fmc_la[8:8] = fmc_la[8:8];
  assign page1_fmc_la[25:25] = fmc_la[25:25];
  assign page1_fmc_la[7:7] = fmc_la[7:7];
  assign page1_fmc_la[4:4] = fmc_la[4:4];
  assign page1_fmc_la[12:12] = fmc_la[12:12];
  assign page1_fmc_la[16:16] = fmc_la[16:16];
  assign page1_fmc_la[20:20] = fmc_la[20:20];
  assign page1_fmc_la[15:15] = fmc_la[15:15];
  assign page1_fmc_la[17:17] = fmc_la[17:17];
  assign page1_fmc_la[23:23] = fmc_la[23:23];
  assign page1_fmc_la[1:1] = fmc_la[1:1];
  assign page1_fmc_la[22:22] = fmc_la[22:22];
  assign page1_fmc_la[11:11] = fmc_la[11:11];
  assign page1_fmc_la[33:0] = fmc_la[33:0];
  assign \page1_fmc_la* [5:5] = \fmc_la* [5:5];
  assign \page1_fmc_la* [17:17] = \fmc_la* [17:17];
  assign \page1_fmc_la* [30:30] = \fmc_la* [30:30];
  assign \page1_fmc_la* [31:31] = \fmc_la* [31:31];
  assign \page1_fmc_la* [29:29] = \fmc_la* [29:29];
  assign \page1_fmc_la* [25:25] = \fmc_la* [25:25];
  assign \page1_fmc_la* [0:0] = \fmc_la* [0:0];
  assign \page1_fmc_la* [6:6] = \fmc_la* [6:6];
  assign \page1_fmc_la* [10:10] = \fmc_la* [10:10];
  assign \page1_fmc_la* [14:14] = \fmc_la* [14:14];
  assign \page1_fmc_la* [18:18] = \fmc_la* [18:18];
  assign \page1_fmc_la* [27:27] = \fmc_la* [27:27];
  assign \page1_fmc_la* [26:26] = \fmc_la* [26:26];
  assign \page1_fmc_la* [24:24] = \fmc_la* [24:24];
  assign \page1_fmc_la* [32:32] = \fmc_la* [32:32];
  assign \page1_fmc_la* [11:11] = \fmc_la* [11:11];
  assign \page1_fmc_la* [21:21] = \fmc_la* [21:21];
  assign \page1_fmc_la* [28:28] = \fmc_la* [28:28];
  assign \page1_fmc_la* [19:19] = \fmc_la* [19:19];
  assign \page1_fmc_la* [22:22] = \fmc_la* [22:22];
  assign \page1_fmc_la* [3:3] = \fmc_la* [3:3];
  assign \page1_fmc_la* [8:8] = \fmc_la* [8:8];
  assign \page1_fmc_la* [12:12] = \fmc_la* [12:12];
  assign \page1_fmc_la* [16:16] = \fmc_la* [16:16];
  assign \page1_fmc_la* [15:15] = \fmc_la* [15:15];
  assign \page1_fmc_la* [23:23] = \fmc_la* [23:23];
  assign \page1_fmc_la* [13:13] = \fmc_la* [13:13];
  assign \page1_fmc_la* [9:9] = \fmc_la* [9:9];
  assign \page1_fmc_la* [1:1] = \fmc_la* [1:1];
  assign \page1_fmc_la* [33:33] = \fmc_la* [33:33];
  assign \page1_fmc_la* [20:20] = \fmc_la* [20:20];
  assign \page1_fmc_la* [7:7] = \fmc_la* [7:7];
  assign \page1_fmc_la* [4:4] = \fmc_la* [4:4];
  assign \page1_fmc_la* [2:2] = \fmc_la* [2:2];
  assign \page1_fmc_la* [33:0] = \fmc_la* [33:0];
  assign page1_fmc_prsnt_m2c_l = fmc_prsnt_m2c_l;
  assign page1_fmc_pwr_good_flash_rst_b = fmc_pwr_good_flash_rst_b;
  assign page1_fmc_tck_buf = fmc_tck_buf;
  assign page1_fmc_tdo = fmc_tdo;
  assign page1_fmc_tms_buf = fmc_tms_buf;
  assign page1_fpga_tdo = fpga_tdo;
  assign page1_ga0 = ga0;
  assign page1_ga1 = ga1;
  assign page1_gbtclk0_m2c = gbtclk0_m2c;
  assign \page1_gbtclk0_m2c*  = \gbtclk0_m2c* ;
  assign page1_gnd = gnd;
  assign page1_iic_scl_main = iic_scl_main;
  assign page1_iic_sda_main = iic_sda_main;
  assign page1_p12v = p12v;
  assign page1_p2v5 = p2v5;
  assign page1_p3v3 = p3v3;
  assign page1_trst_l = trst_l;
  assign page1_vref_a_m2c = vref_a_m2c;

// begin instances 

  con160p_40cdgh page1_i1  (.g({gnd, p2v5, gnd, \fmc_la* [33], fmc_la[33], gnd, \fmc_la* [31], fmc_la[31],
	gnd, \fmc_la* [29], fmc_la[29], gnd, \fmc_la* [25], fmc_la[25], gnd, \fmc_la* [22],
	fmc_la[22], gnd, \fmc_la* [20], fmc_la[20], gnd, \fmc_la* [16], fmc_la[16],
	gnd, \fmc_la* [12], fmc_la[12], gnd, \fmc_la* [8], fmc_la[8], gnd, \fmc_la* [3],
	fmc_la[3], gnd, \fmc_la* [0], fmc_la[0], gnd, gnd, \fmc_clk1_m2c* , fmc_clk1_m2c,
	gnd}),
	.h({p2v5, gnd, \fmc_la* [32], fmc_la[32], gnd, \fmc_la* [30], fmc_la[30],
	gnd, \fmc_la* [28], fmc_la[28], gnd, \fmc_la* [24], fmc_la[24], gnd, \fmc_la* [21],
	fmc_la[21], gnd, \fmc_la* [19], fmc_la[19], gnd, \fmc_la* [15], fmc_la[15],
	gnd, \fmc_la* [11], fmc_la[11], gnd, \fmc_la* [7], fmc_la[7], gnd, \fmc_la* [4],
	fmc_la[4], gnd, \fmc_la* [2], fmc_la[2], gnd, \fmc_clk0_m2c* , fmc_clk0_m2c,
	gnd, fmc_prsnt_m2c_l, vref_a_m2c}),
	.c(/* unconnected */),
	.d(/* unconnected */));

  con160p_40cdgh page1_i2  (.c({gnd, p3v3, gnd, p12v, gnd, p12v, ga0,
	gnd, gnd, iic_sda_main, iic_scl_main, gnd, gnd, \fmc_la* [27], fmc_la[27],
	gnd, gnd, \fmc_la* [18], fmc_la[18], gnd, gnd, \fmc_la* [14], fmc_la[14],
	gnd, gnd, \fmc_la* [10], fmc_la[10], gnd, gnd, \fmc_la* [6], fmc_la[6],
	gnd, gnd, \dp0_m2c* , dp0_m2c, gnd, gnd, \dp0_c2m* , dp0_c2m, gnd}),
	.d({p3v3,
	gnd, p3v3, gnd, p3v3, ga1, trst_l, fmc_tms_buf, p3v3, fmc_tdo, fpga_tdo,
	fmc_tck_buf, gnd, \fmc_la* [26], fmc_la[26], gnd, \fmc_la* [23], fmc_la[23],
	gnd, \fmc_la* [17], fmc_la[17], gnd, \fmc_la* [13], fmc_la[13], gnd, \fmc_la* [9],
	fmc_la[9], gnd, \fmc_la* [5], fmc_la[5], gnd, \fmc_la* [1], fmc_la[1],
	gnd, gnd, \gbtclk0_m2c* , gbtclk0_m2c, gnd, gnd, fmc_pwr_good_flash_rst_b}),
	.g(/* unconnected */),
	.h(/* unconnected */));

endmodule // pc036a_fmc_lpc_connector(sch_1) 
